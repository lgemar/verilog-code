module averager(
	cclk, rstb, ena,
	raw,
	averaged
);

parameter N = 8;
parameter M = 2;

//implement an averager here
// be sure that it only adds to the sum when the ena signal is high

endmodule
